<<<<<<< HEAD
module udp_fulladder(sum,carry,a,b,c);
input a,b,c;
output sum,carry;
udp_sum s1(sum,a,b,c);
udp_carry c1(carry,a,b,c);

=======
module udp_fulladder(sum,carry,a,b,c);
input a,b,c;
output sum,carry;
udp_sum s1(sum,a,b,c);
udp_carry c1(carry,a,b,c);

>>>>>>> d5771bfc649faa2ad63436b77cef34935263306d
endmodule